netcdf small {variables: byte t; data: t = 1;}
