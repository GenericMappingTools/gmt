netcdf bigf2 {
                // fixed-size variables only, large last variable
                // should fail with classic format due to 4 GB var
                // should work fine with 64-bit offset format
dimensions:
	x = 1000 ;
	y = 1000 ;
	z = 1000 ;
variables:
	float x(x) ;
	float y(y) ;
	float z(z) ;
	float fvar(x, y, z) ; // 4 GB variable
	float flast ;
data:
	flast = 42;
}
