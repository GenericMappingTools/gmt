netcdf bigr2 {
                // large last record variable
                // should fail with classic format
                // should work fine with 64-bit offset format
dimensions:
	x = 1000 ;
	y = 1000 ;
	z = 1000 ;
	t = UNLIMITED ;
variables:
	float x(x) ;
	float y(y) ;
	float z(z) ;
	float t(t) ;
	float var2(t, x, y, z) ;  // 4 GB in each record
	float var1(t) ;
data:
	var1 = 42 ;
}
