netcdf ref_tst_opaque_data {
types:
  opaque(10) raw_obs_t ;
  opaque(3) raw_obs2_t ;
dimensions:
	time = 5 ;
variables:
	raw_obs_t raw_obs(time) ;
		raw_obs_t raw_obs:_FillValue = 0XCAFEBABECAFEBABECAF ;
	raw_obs2_t raw_obs2(time) ;
		raw_obs2_t raw_obs2:_FillValue = 0XABC;
data:

 raw_obs = 0X02030405060708090A0B, 0XAABBCCDDEEFFEEDDC, 
    0XFFFFFFFFFFFFFFFFFFFF, _, 0XCF0DEFACED0CAFE0FACA ;
 raw_obs2 = 0X123, _, 0XFFF, _, 0X357 ;
}
