netcdf bigf1 {
                // fixed-size variables only, large last variable
                // should work fine with classic format
                // should work fine with 64-bit offset format
dimensions:
	x = 100 ;
	y = 100 ;
	z = 100 ;
variables:
	float x(x) ;
	float y(y) ;
	float z(z) ;
	float fvar(x, y, z) ;  // 4 GB OK since last fixed-size variable
}
