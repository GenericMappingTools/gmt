netcdf ref_const_test {
dimensions:
  d3=3;
  d4=4;
variables:
    char charv;
    byte int8v(d4);
    short int16v(d3);
    int int32v(d3);
    int64 int64v(d3);
    ubyte uint8v(d4);
    ushort uint16v(d3);
    uint uint32v(d3);
    uint64 uint64v(d3);
    float floatv;
    double doublev;
data:

 charv = 'a';

 int8v = -5b, 5b, 0xaf, 'a';

 int16v = -2000s, 32767s, 0xabcdS;

 int32v = -200000, 256000, 0xabcdabcL;

 int64v = -200000000000L, 51200000000L, 0xabcdabcdabcdabcdL;

 uint8v = -5b, 5b, 0xaf, 'a';

 uint16v = -2000s, 65535s, 0xabcdS;

 uint32v = -200000, 256000, 0xabcdabcL;

 uint64v = -200000000000, 51200000000, 0xabcdabcdabcdabcdL;

 floatv = 516.0f;

 doublev = -77777777.8888;
}
