netcdf test0 {

dimensions:
	i = 2;
	j = 3;
	k = unlimited;
        l = 3 ;

variables:
	char broiled(i,j,l);
		broiled:act = "text string\n\t123";
		broiled:acb = 10b;
		broiled:acs = -200s ;
		broiled:acl = 17000 ;
		broiled:acf = -2.0f, 1.f, 0.0f ;
		broiled:acd = -1.0, 2.7182818284590455;
	byte the_bullet(i,j);
	short order(i,j);
	int rigue(i,j);
	float a_loan(i,j);
	double entendre(i,j);
	char cscalar;
	double dscalar;
	char cnodata(i);
	byte bnodata(i);
	short snodata(i);
	int inodata(i);
	float fnodata(i);
	double dnodata(i);
	int i(i);
	float j(j);
	byte l(l);

	:glob = "Global attribute" ;

data:
	broiled = "indistinguishable" ;
	the_bullet = -127,0,127,128,255;
	order = 1s, 2s, 3s, 4s, 5s, 6s;
	rigue = 2, 3, 4, 5, 6, 7 ;
	a_loan = 3.f, 4.f, 5.f, 6.f, 7.f, 1.0e12f ;
	entendre = '\4', 5s, 6, 7.0f, 8.0, 1.0e30 ;
	i = 10, 20;
	j = 2, 4, 6;
	l = 10, 9, 8;
}
