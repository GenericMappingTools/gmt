netcdf nc_sync {
    dimensions:
	dim0 = 53;
	dim1 = 67;
	dim2 = 30;
	dim3 = UNLIMITED ; // (0 currently)
    variables:
	double var0(dim3,dim2,dim1,dim0);
	double var1(dim3,dim2,dim1,dim0);
	double var2(dim3,dim2,dim1,dim0);
	double var3(dim3,dim2,dim1,dim0);
	double var4(dim3,dim2,dim1,dim0);
	double var5(dim3,dim2,dim1,dim0);
	double var6(dim3,dim2,dim1,dim0);
	double var7(dim3,dim2,dim1,dim0);
	double var8(dim3,dim2,dim1,dim0);
	double var9(dim3,dim2,dim1,dim0);
	double var10(dim3,dim2,dim1,dim0);
	double var11(dim3,dim2,dim1,dim0);
	double var12(dim3,dim2,dim1,dim0);
	double var13(dim3,dim2,dim1,dim0);
	double var14(dim3,dim2,dim1,dim0);
	double var15(dim3,dim2,dim1,dim0);
	double var16(dim3,dim2,dim1,dim0);
	double var17(dim3,dim2,dim1,dim0);
	double var18(dim3,dim2,dim1,dim0);
	double var19(dim3,dim2,dim1,dim0);
	double var20(dim3,dim2,dim1,dim0);
	double var21(dim3,dim2,dim1,dim0);
	double var22(dim3,dim2,dim1,dim0);
	double var23(dim3,dim2,dim1,dim0);
	double var24(dim3,dim2,dim1,dim0);
	double var25(dim3,dim2,dim1,dim0);
	double var26(dim3,dim2,dim1,dim0);
	double var27(dim3,dim2,dim1,dim0);
	double var28(dim3,dim2,dim1,dim0);
	double var29(dim3,dim2,dim1,dim0);
	double var30(dim3,dim2,dim1,dim0);
	double var31(dim3,dim2,dim1,dim0);
	double var32(dim3,dim2,dim1,dim0);
	double var33(dim3,dim2,dim1,dim0);
	double var34(dim3,dim2,dim1,dim0);
	double var35(dim3,dim2,dim1,dim0);
	double var36(dim3,dim2,dim1,dim0);
data:
}
