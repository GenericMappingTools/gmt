netcdf ref_tst_compounds3 {
types:
  compound cmp_t {
    float x ;
    double y ;
  }; // cmp_t
dimensions:
	n = 1 ;
variables:
	cmp_t var(n) ;
data:

 var = {1, -2} ;
}
