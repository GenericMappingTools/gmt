netcdf ref_tst_small {
dimensions:
	Time = UNLIMITED ; // (2 currently)
	DateStrLen = 19 ;
variables:
	char Times(Time, DateStrLen) ;

// global attributes:
		:TITLE = " OUTPUT FROM WRF V2.0.3.1 MODEL" ;
data:

 Times =
  "2005-04-11_12:00:00",
  "2005-04-11_13:00:00" ;
}
