netcdf ref_nctst_64bit_offset {
dimensions:
	lat = 4 ;
	lon = 3 ;
	frtime = UNLIMITED ; // (2 currently)
	timelen = 20 ;
variables:
	float P(frtime, lat, lon) ;
		P:long_name = "pressure at maximum wind" ;
		P:units = "hectopascals" ;
		P:valid_range = 0.f, 1500.f ;
		P:_FillValue = -9999.f ;
	float lat(lat) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
	float lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
	int frtime(frtime) ;
		frtime:long_name = "forecast time" ;
		frtime:units = "hours" ;
	char reftime(timelen) ;
		reftime:long_name = "reference time" ;
		reftime:units = "text_time" ;
	int scalarv ;
		scalarv:scalar_att = 1 ;

// global attributes:
		:history = "created by Unidata LDM from NPS broadcast" ;
		:title = "NMC Global Product Set: Pressure at Maximum Wind" ;
data:

 P =
  950, 951, 952,
  953, 954, 955,
  956, 957, 958,
  959, 960, 961,
  962, 963, 964,
  965, 966, 967,
  968, 969, 970,
  971, 972, 973 ;

 lat = -90, -87.5, -85, -82.5 ;

 lon = -180, -175, -170 ;

 frtime = 12, 18 ;

 reftime = "1992-3-21 12:00" ;

 scalarv = _ ;
}
