netcdf tst_ncml {
dimensions:
   m = 2;
   t = unlimited;
variables:
   float var (t, m);
     var:tatt = "text attribute value" ;
     var:natt = 1, 2;
   :gtatt = "<, >, \', \", and &" ;
   :gnatt = 3, 4;
}
