netcdf fills {
dimensions:
	n = 2 ;
variables:
	double d(n) ;
	float f(n) ;
	int l(n) ;
	short s(n) ;
	byte b(n) ;
data:

 d = 1, _ ;

 f = 1, _ ;

 l = 1, _ ;

 s = 1, _ ;

 b = 1, -127 ;
}
