netcdf tst_comp2 {
types:
  compound vecmat_t {
    char day ;
    char mnth(3) ;
    short vect(3) ;
    float matr(2, 3) ;
  }; // vecmat_t
dimensions:
	n = 3 ;
variables:
	vecmat_t obs(n) ;
		vecmat_t obs:_FillValue = {"?", {"---"}, {-1, -2, -3}, {-4, -5, -6, -7, -8, -9}} ;
data:

 obs = {"S", {"jan"}, {1, 2, 3}, {4, 5, 6, 7, 8, 9}}, 
    {"M", {"feb"}, {11, 12, 13}, {4.25, 5.25, 6.25, 7.25, 8.25, 9.25}}, 
    {"T", {"mar"}, {21, 22, 23}, {4.5, 5.5, 6.5, 7.5, 8.5, 9.5}} ;
}
