netcdf small2 {
dimensions:
	t = UNLIMITED ;
	m = 5 ;
variables:
	byte b(t, m) ;
data:

 b = 1, 2, 3, 4, 5 ;
}
