netcdf ref_tst_vlen_data { // H/T to Lynton Appel for extra tests of vlen
types:
  float(*) row_of_floats ;
  int(*) vlen_int ;
  compound singleCompoundType {
    vlen_int vlenIntVector(2) ;
  }; // singleCompoundType
  compound pfCoilType {
    vlen_int name ;
  }; // pfCoilType
  pfCoilType(*) vlen_t ;
  vlen_int(*) vlen_int2 ;
  compound singleCompoundType2 {
    vlen_int2 vlenIntVector ;
  }; // singleCompoundType2
dimensions:
	m = 5 ;
	vlenDim = 2 ;
variables:
	row_of_floats ragged_array(m) ;
		row_of_floats ragged_array:_FillValue = {-999} ;
	vlen_int vdata ;
	singleCompoundType singleCompound ;
	vlen_t pfCircuits ;
	singleCompoundType2 singleCompound2 ;
	vlen_int vlenIntVector(vlenDim) ;
data:

 ragged_array = {10, 11, 12, 13, 14}, {20, 21, 22, 23}, {30, 31, 32}, 
    {40, 41}, _ ;

 vdata = {1, 2, 3} ;

 singleCompound = {{{11}, {12}}} ;

 pfCircuits = {{{1, 2, 3}}, {{2}}, {{3}}, {{4}}} ;

 singleCompound2 = {{{11}, {12}}} ;

 vlenIntVector = {1, 2, 3}, {1, 2, 3} ;
}
