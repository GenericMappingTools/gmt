netcdf bigf1 {
                // fixed-size variables only, large last variable
                // should work fine with classic format
                // should work fine with 64-bit offset format
dimensions:
	x = 1000 ;
	y = 1000 ;
	z = 1000 ;
variables:
	float x(x) ;
	float y(y) ;
	float z(z) ;
	float fvar(x, y, z) ;  // 4 GB OK since last fixed-size variable
}
