netcdf ref_tst_unlim2 {
dimensions:
  D2  = 2 ;
  U1  = UNLIMITED ; // (1 currently)
  U2  = UNLIMITED ; // (2 currently)
  UU3 = UNLIMITED ; // (4 currently)
  UUU2 = UNLIMITED ; // (2 currently)
  UUU3 = UNLIMITED ; // (6 currently)
variables:
  char cuu(U1,D2,UU3);
  char cuuu(U2,UUU2,UUU3);
data:
  cuu  = {"a","def"},{"xy"} ;
  cuuu = {{"1", "two"}}, {{"three"},{"four","xy"}} ;
}


