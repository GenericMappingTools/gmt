netcdf tst_opaque_data {
types:
  opaque(11) raw_obs_t ;
dimensions:
	time = 5 ;
variables:
	raw_obs_t raw_obs(time) ;
		raw_obs_t raw_obs:_FillValue = 0XCAFEBABECAFEBABECAFEBA ;
data:

 raw_obs = 0X0102030405060708090A0B, 0XAABBCCDDEEFFEEDDCCBBAA, 
    0XFFFFFFFFFFFFFFFFFFFFFF, _, 0XCF0DEFACED0CAFE0FACADE ;
}
