netcdf ref_tst_group_data {
dimensions:
	dim = 4 ;
variables:
	float var(dim) ;
		var:units = "m/s" ;

// global attributes:
		:title = "for testing groups" ;
data:

 var = 1, 2, 3, 4 ;

group: g1 {
  dimensions:
  	dim = 1 ;
  variables:
  	float var(dim) ;
  		var:units = "km/hour" ;

  // global attributes:
  		:title = "in first group" ;
  data:

   var = 1 ;
  } // group g1

group: g2 {
  dimensions:
  	dim = 2 ;
  variables:
  	float var(dim) ;
  		var:units = "cm/sec" ;

  // global attributes:
  		:title = "in second group" ;
  data:

   var = 1, 2 ;

  group: g3 {
    dimensions:
    	dim = 3 ;
    variables:
    	float var(dim) ;
    		var:units = "mm/msec" ;

    // global attributes:
    		:title = "in third group" ;
    data:

     var = 1, 2, 3 ;
    } // group g3
  } // group g2
}
