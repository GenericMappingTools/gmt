netcdf tst_nans {
dimensions:
	dim = 3 ;
variables:
	float fvar(dim) ;
		fvar:_FillValue = NaNf ;
		fvar:att = -Infinityf, NaNf, Infinityf ;
	double dvar(dim) ;
		dvar:_FillValue = NaN ;
		dvar:att = -Infinity, NaN, Infinity ;
data:

 fvar = -Infinityf, _, Infinityf ;

 dvar = -Infinity, _, Infinity ;
}
