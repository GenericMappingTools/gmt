netcdf tst_chunks {
dimensions:
	dim1 = 6 ;
	dim2 = 12 ;
	dim3 = 4 ;
variables:
	float var_contiguous(dim1, dim2, dim3) ;
		var_contiguous:_Storage = "contiguous" ;
	float var_chunked(dim1, dim2, dim3) ;
		var_chunked:_Storage = "chunked" ;
		var_chunked:_ChunkSizes = 2, 3, 1 ;
	float var_compressed(dim1, dim2, dim3) ;
		var_compressed:_Storage = "chunked" ;
		var_compressed:_ChunkSizes = 2, 3, 1 ;
		var_compressed:_DeflateLevel = 1 ;

// global attributes:
		:_Format = "netCDF-4 classic model" ;
data:

 var_contiguous =
  0, 0, 0, 0,
  1, 1, 1, 1,
  2, 2, 2, 2,
  3, 3, 3, 3,
  4, 4, 4, 4,
  5, 5, 5, 5,
  6, 6, 6, 6,
  7, 7, 7, 7,
  8, 8, 8, 8,
  9, 9, 9, 9,
  10, 10, 10, 10,
  11, 11, 11, 11,
  12, 12, 12, 12,
  13, 13, 13, 13,
  14, 14, 14, 14,
  15, 15, 15, 15,
  16, 16, 16, 16,
  17, 17, 17, 17,
  18, 18, 18, 18,
  19, 19, 19, 19,
  20, 20, 20, 20,
  21, 21, 21, 21,
  22, 22, 22, 22,
  23, 23, 23, 23,
  24, 24, 24, 24,
  25, 25, 25, 25,
  26, 26, 26, 26,
  27, 27, 27, 27,
  28, 28, 28, 28,
  29, 29, 29, 29,
  30, 30, 30, 30,
  31, 31, 31, 31,
  32, 32, 32, 32,
  33, 33, 33, 33,
  34, 34, 34, 34,
  35, 35, 35, 35,
  36, 36, 36, 36,
  37, 37, 37, 37,
  38, 38, 38, 38,
  39, 39, 39, 39,
  40, 40, 40, 40,
  41, 41, 41, 41,
  42, 42, 42, 42,
  43, 43, 43, 43,
  44, 44, 44, 44,
  45, 45, 45, 45,
  46, 46, 46, 46,
  47, 47, 47, 47,
  48, 48, 48, 48,
  49, 49, 49, 49,
  50, 50, 50, 50,
  51, 51, 51, 51,
  52, 52, 52, 52,
  53, 53, 53, 53,
  54, 54, 54, 54,
  55, 55, 55, 55,
  56, 56, 56, 56,
  57, 57, 57, 57,
  58, 58, 58, 58,
  59, 59, 59, 59,
  60, 60, 60, 60,
  61, 61, 61, 61,
  62, 62, 62, 62,
  63, 63, 63, 63,
  64, 64, 64, 64,
  65, 65, 65, 65,
  66, 66, 66, 66,
  67, 67, 67, 67,
  68, 68, 68, 68,
  69, 69, 69, 69,
  70, 70, 70, 70,
  71, 71, 71, 71 ;

 var_chunked =
  0, 0, 0, 0,
  1, 1, 1, 1,
  2, 2, 2, 2,
  3, 3, 3, 3,
  4, 4, 4, 4,
  5, 5, 5, 5,
  6, 6, 6, 6,
  7, 7, 7, 7,
  8, 8, 8, 8,
  9, 9, 9, 9,
  10, 10, 10, 10,
  11, 11, 11, 11,
  12, 12, 12, 12,
  13, 13, 13, 13,
  14, 14, 14, 14,
  15, 15, 15, 15,
  16, 16, 16, 16,
  17, 17, 17, 17,
  18, 18, 18, 18,
  19, 19, 19, 19,
  20, 20, 20, 20,
  21, 21, 21, 21,
  22, 22, 22, 22,
  23, 23, 23, 23,
  24, 24, 24, 24,
  25, 25, 25, 25,
  26, 26, 26, 26,
  27, 27, 27, 27,
  28, 28, 28, 28,
  29, 29, 29, 29,
  30, 30, 30, 30,
  31, 31, 31, 31,
  32, 32, 32, 32,
  33, 33, 33, 33,
  34, 34, 34, 34,
  35, 35, 35, 35,
  36, 36, 36, 36,
  37, 37, 37, 37,
  38, 38, 38, 38,
  39, 39, 39, 39,
  40, 40, 40, 40,
  41, 41, 41, 41,
  42, 42, 42, 42,
  43, 43, 43, 43,
  44, 44, 44, 44,
  45, 45, 45, 45,
  46, 46, 46, 46,
  47, 47, 47, 47,
  48, 48, 48, 48,
  49, 49, 49, 49,
  50, 50, 50, 50,
  51, 51, 51, 51,
  52, 52, 52, 52,
  53, 53, 53, 53,
  54, 54, 54, 54,
  55, 55, 55, 55,
  56, 56, 56, 56,
  57, 57, 57, 57,
  58, 58, 58, 58,
  59, 59, 59, 59,
  60, 60, 60, 60,
  61, 61, 61, 61,
  62, 62, 62, 62,
  63, 63, 63, 63,
  64, 64, 64, 64,
  65, 65, 65, 65,
  66, 66, 66, 66,
  67, 67, 67, 67,
  68, 68, 68, 68,
  69, 69, 69, 69,
  70, 70, 70, 70,
  71, 71, 71, 71 ;

 var_compressed =
  0, 0, 0, 0,
  1, 1, 1, 1,
  2, 2, 2, 2,
  3, 3, 3, 3,
  4, 4, 4, 4,
  5, 5, 5, 5,
  6, 6, 6, 6,
  7, 7, 7, 7,
  8, 8, 8, 8,
  9, 9, 9, 9,
  10, 10, 10, 10,
  11, 11, 11, 11,
  12, 12, 12, 12,
  13, 13, 13, 13,
  14, 14, 14, 14,
  15, 15, 15, 15,
  16, 16, 16, 16,
  17, 17, 17, 17,
  18, 18, 18, 18,
  19, 19, 19, 19,
  20, 20, 20, 20,
  21, 21, 21, 21,
  22, 22, 22, 22,
  23, 23, 23, 23,
  24, 24, 24, 24,
  25, 25, 25, 25,
  26, 26, 26, 26,
  27, 27, 27, 27,
  28, 28, 28, 28,
  29, 29, 29, 29,
  30, 30, 30, 30,
  31, 31, 31, 31,
  32, 32, 32, 32,
  33, 33, 33, 33,
  34, 34, 34, 34,
  35, 35, 35, 35,
  36, 36, 36, 36,
  37, 37, 37, 37,
  38, 38, 38, 38,
  39, 39, 39, 39,
  40, 40, 40, 40,
  41, 41, 41, 41,
  42, 42, 42, 42,
  43, 43, 43, 43,
  44, 44, 44, 44,
  45, 45, 45, 45,
  46, 46, 46, 46,
  47, 47, 47, 47,
  48, 48, 48, 48,
  49, 49, 49, 49,
  50, 50, 50, 50,
  51, 51, 51, 51,
  52, 52, 52, 52,
  53, 53, 53, 53,
  54, 54, 54, 54,
  55, 55, 55, 55,
  56, 56, 56, 56,
  57, 57, 57, 57,
  58, 58, 58, 58,
  59, 59, 59, 59,
  60, 60, 60, 60,
  61, 61, 61, 61,
  62, 62, 62, 62,
  63, 63, 63, 63,
  64, 64, 64, 64,
  65, 65, 65, 65,
  66, 66, 66, 66,
  67, 67, 67, 67,
  68, 68, 68, 68,
  69, 69, 69, 69,
  70, 70, 70, 70,
  71, 71, 71, 71 ;
}
