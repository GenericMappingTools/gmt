netcdf nc_test_netcdf4 {
dimensions:
	Dr = UNLIMITED ; // (2 currently)
	D1 = 1 ;
	D2 = 2 ;
	D3 = 3 ;
	D4 = 4 ;
variables:
	char c ;
	byte b ;
		b:c = "" ;
	short s ;
		s:b = -128b ;
		s:s = -32768s, 32767s ;
	int i ;
		i:i = -2147483648, 2147483647, -2147483648 ;
		i:f = -3.402823e+38f, 3.402823e+38f, -Infinityf, Infinityf ;
		i:d = -1.79769313486232e+308, 1.79769313486232e+308, -1., 1., 660. ;
	float f ;
	double d ;
		d:c = "�\177AZ$&" ;
	char cr(Dr) ;
	byte br(Dr) ;
	short sr(Dr) ;
	int ir(Dr) ;
	float fr(Dr) ;
	double dr(Dr) ;
	char c1(D1) ;
	byte b1(D1) ;
	short s1(D1) ;
	int i1(D1) ;
	float f1(D1) ;
	double d1(D1) ;
	char c2(D2) ;
	byte b2(D2) ;
	short s2(D2) ;
	int i2(D2) ;
	float f2(D2) ;
	double d2(D2) ;
	char c3(D3) ;
	byte b3(D3) ;
	short s3(D3) ;
	int i3(D3) ;
	float f3(D3) ;
	double d3(D3) ;
	char c4(D4) ;
	byte b4(D4) ;
	short s4(D4) ;
	int i4(D4) ;
	float f4(D4) ;
	double d4(D4) ;
	char cr1(Dr, D1) ;
	byte br2(Dr, D2) ;
	short sr3(Dr, D3) ;
	int ir4(Dr, D4) ;
	float f11(D1, D1) ;
	double d12(D1, D2) ;
	char c13(D1, D3) ;
	byte b14(D1, D4) ;
	short s21(D2, D1) ;
	int i22(D2, D2) ;
	float f23(D2, D3) ;
	double d24(D2, D4) ;
	char c31(D3, D1) ;
	byte b32(D3, D2) ;
	short s33(D3, D3) ;
	int i34(D3, D4) ;
	float f41(D4, D1) ;
	double d42(D4, D2) ;
	char c43(D4, D3) ;
	byte b44(D4, D4) ;
	short sr11(Dr, D1, D1) ;
	int ir12(Dr, D1, D2) ;
	float fr13(Dr, D1, D3) ;
	double dr14(Dr, D1, D4) ;
	char cr21(Dr, D2, D1) ;
	byte br22(Dr, D2, D2) ;
	short sr23(Dr, D2, D3) ;
	int ir24(Dr, D2, D4) ;
	float fr31(Dr, D3, D1) ;
	double dr32(Dr, D3, D2) ;
	char cr33(Dr, D3, D3) ;
	byte br34(Dr, D3, D4) ;
	short sr41(Dr, D4, D1) ;
	int ir42(Dr, D4, D2) ;
	float fr43(Dr, D4, D3) ;
	double dr44(Dr, D4, D4) ;
	char c111(D1, D1, D1) ;
	byte b112(D1, D1, D2) ;
	short s113(D1, D1, D3) ;
	int i114(D1, D1, D4) ;
	float f121(D1, D2, D1) ;
	double d122(D1, D2, D2) ;
	char c123(D1, D2, D3) ;
	byte b124(D1, D2, D4) ;
	short s131(D1, D3, D1) ;
	int i132(D1, D3, D2) ;
	float f133(D1, D3, D3) ;
	double d134(D1, D3, D4) ;
	char c141(D1, D4, D1) ;
	byte b142(D1, D4, D2) ;
	short s143(D1, D4, D3) ;
	int i144(D1, D4, D4) ;
	float f211(D2, D1, D1) ;
	double d212(D2, D1, D2) ;
	char c213(D2, D1, D3) ;
	byte b214(D2, D1, D4) ;
	short s221(D2, D2, D1) ;
	int i222(D2, D2, D2) ;
	float f223(D2, D2, D3) ;
	double d224(D2, D2, D4) ;
	char c231(D2, D3, D1) ;
	byte b232(D2, D3, D2) ;
	short s233(D2, D3, D3) ;
	int i234(D2, D3, D4) ;
	float f241(D2, D4, D1) ;
	double d242(D2, D4, D2) ;
	char c243(D2, D4, D3) ;
	byte b244(D2, D4, D4) ;
	short s311(D3, D1, D1) ;
	int i312(D3, D1, D2) ;
	float f313(D3, D1, D3) ;
	double d314(D3, D1, D4) ;
	char c321(D3, D2, D1) ;
	byte b322(D3, D2, D2) ;
	short s323(D3, D2, D3) ;
	int i324(D3, D2, D4) ;
	float f331(D3, D3, D1) ;
	double d332(D3, D3, D2) ;
	char c333(D3, D3, D3) ;
	byte b334(D3, D3, D4) ;
	short s341(D3, D4, D1) ;
	int i342(D3, D4, D2) ;
	float f343(D3, D4, D3) ;
	double d344(D3, D4, D4) ;
	char c411(D4, D1, D1) ;
	byte b412(D4, D1, D2) ;
	short s413(D4, D1, D3) ;
	int i414(D4, D1, D4) ;
	float f421(D4, D2, D1) ;
	double d422(D4, D2, D2) ;
	char c423(D4, D2, D3) ;
	byte b424(D4, D2, D4) ;
	short s431(D4, D3, D1) ;
	int i432(D4, D3, D2) ;
	float f433(D4, D3, D3) ;
	double d434(D4, D3, D4) ;
	char c441(D4, D4, D1) ;
	byte b442(D4, D4, D2) ;
	short s443(D4, D4, D3) ;
	int i444(D4, D4, D4) ;

// global attributes:
		:Gc = "�" ;
		:Gb = -128b, 127b ;
		:Gs = -32768s, 32767s, 32767s ;
		:Gi = -2147483648, 2147483647, -2147483648, -2147483648 ;
		:Gf = -3.402823e+38f, 3.402823e+38f, -Infinityf, Infinityf, 531.f ;
		:Gd = -1.79769313486232e+308, 1.79769313486232e+308, -1., 1., 660., 650. ;
data:

 c = "\002" ;

 b = -2 ;

 s = -5 ;

 i = -20 ;

 f = -9 ;

 d = -10 ;

 cr = "\200\177" ;

 br = -128, 127 ;

 sr = -32768, 32767 ;

 ir = -2147483648, 2147483647 ;

 fr = -3.402823e+38, 3.402823e+38 ;

 dr = -1.79769313486232e+308, 1.79769313486232e+308 ;

 c1 = "\200" ;

 b1 = -128 ;

 s1 = -32768 ;

 i1 = -2147483648 ;

 f1 = -3.402823e+38 ;

 d1 = -1.79769313486232e+308 ;

 c2 = "\200\177" ;

 b2 = -128, 127 ;

 s2 = -32768, 32767 ;

 i2 = -2147483648, 2147483647 ;

 f2 = -3.402823e+38, 3.402823e+38 ;

 d2 = -1.79769313486232e+308, 1.79769313486232e+308 ;

 c3 = "\200\177A" ;

 b3 = -128, 127, 127 ;

 s3 = -32768, 32767, 32767 ;

 i3 = -2147483648, 2147483647, -2147483648 ;

 f3 = -3.402823e+38, 3.402823e+38, -Infinityf ;

 d3 = -1.79769313486232e+308, 1.79769313486232e+308, -1 ;

 c4 = "\200\177AZ" ;

 b4 = -128, 127, 127, -128 ;

 s4 = -32768, 32767, 32767, -32768 ;

 i4 = -2147483648, 2147483647, -2147483648, -2147483648 ;

 f4 = -3.402823e+38, 3.402823e+38, -Infinityf, Infinityf ;

 d4 = -1.79769313486232e+308, 1.79769313486232e+308, -1, 1 ;

 cr1 =
  "\030",
  "\034" ;

 br2 =
  -24, -26,
  -20, -22 ;

 sr3 =
  -375, -380, -385,
  -350, -355, -360 ;

 ir4 =
  -24000, -24020, -24040, -24060,
  -23600, -23620, -23640, -23660 ;

 f11 =
  -2187 ;

 d12 =
  -3000, -3010 ;

 c13 =
  "\030\032\034" ;

 b14 =
  -24, -26, -28, -30 ;

 s21 =
  -375,
  -350 ;

 i22 =
  -24000, -24020,
  -23600, -23620 ;

 f23 =
  -2187, -2196, -2205,
  -2106, -2115, -2124 ;

 d24 =
  -3000, -3010, -3020, -3030,
  -2900, -2910, -2920, -2930 ;

 c31 =
  "\030",
  "\034",
  " " ;

 b32 =
  -24, -26,
  -20, -22,
  -16, -18 ;

 s33 =
  -375, -380, -385,
  -350, -355, -360,
  -325, -330, -335 ;

 i34 =
  -24000, -24020, -24040, -24060,
  -23600, -23620, -23640, -23660,
  -23200, -23220, -23240, -23260 ;

 f41 =
  -2187,
  -2106,
  -2025,
  -1944 ;

 d42 =
  -3000, -3010,
  -2900, -2910,
  -2800, -2810,
  -2700, -2710 ;

 c43 =
  "\030\032\034",
  "\034\036 ",
  " \"$",
  "$&(" ;

 b44 =
  -24, -26, -28, -30,
  -20, -22, -24, -26,
  -16, -18, -20, -22,
  -12, -14, -16, -18 ;

 sr11 =
  2500,
  2375 ;

 ir12 =
  640000, 639980,
  632000, 631980 ;

 fr13 =
  26244, 26235, 26226,
  25515, 25506, 25497 ;

 dr14 =
  40000, 39990, 39980, 39970,
  39000, 38990, 38980, 38970 ;

 cr21 =
  "@",
  "D",
  "H",
  "L" ;

 br22 =
  64, 62,
  68, 66,
  56, 54,
  60, 58 ;

 sr23 =
  2500, 2495, 2490,
  2525, 2520, 2515,
  2375, 2370, 2365,
  2400, 2395, 2390 ;

 ir24 =
  640000, 639980, 639960, 639940,
  640400, 640380, 640360, 640340,
  632000, 631980, 631960, 631940,
  632400, 632380, 632360, 632340 ;

 fr31 =
  26244,
  26325,
  26406,
  25515,
  25596,
  25677 ;

 dr32 =
  40000, 39990,
  40100, 40090,
  40200, 40190,
  39000, 38990,
  39100, 39090,
  39200, 39190 ;

 cr33 =
  "@BD",
  "DFH",
  "HJL",
  "HJL",
  "LNP",
  "PRT" ;

 br34 =
  64, 62, 60, 58,
  68, 66, 64, 62,
  72, 70, 68, 66,
  56, 54, 52, 50,
  60, 58, 56, 54,
  64, 62, 60, 58 ;

 sr41 =
  2500,
  2525,
  2550,
  2575,
  2375,
  2400,
  2425,
  2450 ;

 ir42 =
  640000, 639980,
  640400, 640380,
  640800, 640780,
  641200, 641180,
  632000, 631980,
  632400, 632380,
  632800, 632780,
  633200, 633180 ;

 fr43 =
  26244, 26235, 26226,
  26325, 26316, 26307,
  26406, 26397, 26388,
  26487, 26478, 26469,
  25515, 25506, 25497,
  25596, 25587, 25578,
  25677, 25668, 25659,
  25758, 25749, 25740 ;

 dr44 =
  40000, 39990, 39980, 39970,
  40100, 40090, 40080, 40070,
  40200, 40190, 40180, 40170,
  40300, 40290, 40280, 40270,
  39000, 38990, 38980, 38970,
  39100, 39090, 39080, 39070,
  39200, 39190, 39180, 39170,
  39300, 39290, 39280, 39270 ;

 c111 =
  "@" ;

 b112 =
  64, 62 ;

 s113 =
  2500, 2495, 2490 ;

 i114 =
  640000, 639980, 639960, 639940 ;

 f121 =
  26244,
  26325 ;

 d122 =
  40000, 39990,
  40100, 40090 ;

 c123 =
  "@BD",
  "DFH" ;

 b124 =
  64, 62, 60, 58,
  68, 66, 64, 62 ;

 s131 =
  2500,
  2525,
  2550 ;

 i132 =
  640000, 639980,
  640400, 640380,
  640800, 640780 ;

 f133 =
  26244, 26235, 26226,
  26325, 26316, 26307,
  26406, 26397, 26388 ;

 d134 =
  40000, 39990, 39980, 39970,
  40100, 40090, 40080, 40070,
  40200, 40190, 40180, 40170 ;

 c141 =
  "@",
  "D",
  "H",
  "L" ;

 b142 =
  64, 62,
  68, 66,
  72, 70,
  76, 74 ;

 s143 =
  2500, 2495, 2490,
  2525, 2520, 2515,
  2550, 2545, 2540,
  2575, 2570, 2565 ;

 i144 =
  640000, 639980, 639960, 639940,
  640400, 640380, 640360, 640340,
  640800, 640780, 640760, 640740,
  641200, 641180, 641160, 641140 ;

 f211 =
  26244,
  25515 ;

 d212 =
  40000, 39990,
  39000, 38990 ;

 c213 =
  "@BD",
  "HJL" ;

 b214 =
  64, 62, 60, 58,
  56, 54, 52, 50 ;

 s221 =
  2500,
  2525,
  2375,
  2400 ;

 i222 =
  640000, 639980,
  640400, 640380,
  632000, 631980,
  632400, 632380 ;

 f223 =
  26244, 26235, 26226,
  26325, 26316, 26307,
  25515, 25506, 25497,
  25596, 25587, 25578 ;

 d224 =
  40000, 39990, 39980, 39970,
  40100, 40090, 40080, 40070,
  39000, 38990, 38980, 38970,
  39100, 39090, 39080, 39070 ;

 c231 =
  "@",
  "D",
  "H",
  "H",
  "L",
  "P" ;

 b232 =
  64, 62,
  68, 66,
  72, 70,
  56, 54,
  60, 58,
  64, 62 ;

 s233 =
  2500, 2495, 2490,
  2525, 2520, 2515,
  2550, 2545, 2540,
  2375, 2370, 2365,
  2400, 2395, 2390,
  2425, 2420, 2415 ;

 i234 =
  640000, 639980, 639960, 639940,
  640400, 640380, 640360, 640340,
  640800, 640780, 640760, 640740,
  632000, 631980, 631960, 631940,
  632400, 632380, 632360, 632340,
  632800, 632780, 632760, 632740 ;

 f241 =
  26244,
  26325,
  26406,
  26487,
  25515,
  25596,
  25677,
  25758 ;

 d242 =
  40000, 39990,
  40100, 40090,
  40200, 40190,
  40300, 40290,
  39000, 38990,
  39100, 39090,
  39200, 39190,
  39300, 39290 ;

 c243 =
  "@BD",
  "DFH",
  "HJL",
  "LNP",
  "HJL",
  "LNP",
  "PRT",
  "TVX" ;

 b244 =
  64, 62, 60, 58,
  68, 66, 64, 62,
  72, 70, 68, 66,
  76, 74, 72, 70,
  56, 54, 52, 50,
  60, 58, 56, 54,
  64, 62, 60, 58,
  68, 66, 64, 62 ;

 s311 =
  2500,
  2375,
  2250 ;

 i312 =
  640000, 639980,
  632000, 631980,
  624000, 623980 ;

 f313 =
  26244, 26235, 26226,
  25515, 25506, 25497,
  24786, 24777, 24768 ;

 d314 =
  40000, 39990, 39980, 39970,
  39000, 38990, 38980, 38970,
  38000, 37990, 37980, 37970 ;

 c321 =
  "@",
  "D",
  "H",
  "L",
  "P",
  "T" ;

 b322 =
  64, 62,
  68, 66,
  56, 54,
  60, 58,
  48, 46,
  52, 50 ;

 s323 =
  2500, 2495, 2490,
  2525, 2520, 2515,
  2375, 2370, 2365,
  2400, 2395, 2390,
  2250, 2245, 2240,
  2275, 2270, 2265 ;

 i324 =
  640000, 639980, 639960, 639940,
  640400, 640380, 640360, 640340,
  632000, 631980, 631960, 631940,
  632400, 632380, 632360, 632340,
  624000, 623980, 623960, 623940,
  624400, 624380, 624360, 624340 ;

 f331 =
  26244,
  26325,
  26406,
  25515,
  25596,
  25677,
  24786,
  24867,
  24948 ;

 d332 =
  40000, 39990,
  40100, 40090,
  40200, 40190,
  39000, 38990,
  39100, 39090,
  39200, 39190,
  38000, 37990,
  38100, 38090,
  38200, 38190 ;

 c333 =
  "@BD",
  "DFH",
  "HJL",
  "HJL",
  "LNP",
  "PRT",
  "PRT",
  "TVX",
  "XZ\\" ;

 b334 =
  64, 62, 60, 58,
  68, 66, 64, 62,
  72, 70, 68, 66,
  56, 54, 52, 50,
  60, 58, 56, 54,
  64, 62, 60, 58,
  48, 46, 44, 42,
  52, 50, 48, 46,
  56, 54, 52, 50 ;

 s341 =
  2500,
  2525,
  2550,
  2575,
  2375,
  2400,
  2425,
  2450,
  2250,
  2275,
  2300,
  2325 ;

 i342 =
  640000, 639980,
  640400, 640380,
  640800, 640780,
  641200, 641180,
  632000, 631980,
  632400, 632380,
  632800, 632780,
  633200, 633180,
  624000, 623980,
  624400, 624380,
  624800, 624780,
  625200, 625180 ;

 f343 =
  26244, 26235, 26226,
  26325, 26316, 26307,
  26406, 26397, 26388,
  26487, 26478, 26469,
  25515, 25506, 25497,
  25596, 25587, 25578,
  25677, 25668, 25659,
  25758, 25749, 25740,
  24786, 24777, 24768,
  24867, 24858, 24849,
  24948, 24939, 24930,
  25029, 25020, 25011 ;

 d344 =
  40000, 39990, 39980, 39970,
  40100, 40090, 40080, 40070,
  40200, 40190, 40180, 40170,
  40300, 40290, 40280, 40270,
  39000, 38990, 38980, 38970,
  39100, 39090, 39080, 39070,
  39200, 39190, 39180, 39170,
  39300, 39290, 39280, 39270,
  38000, 37990, 37980, 37970,
  38100, 38090, 38080, 38070,
  38200, 38190, 38180, 38170,
  38300, 38290, 38280, 38270 ;

 c411 =
  "@",
  "H",
  "P",
  "X" ;

 b412 =
  64, 62,
  56, 54,
  48, 46,
  40, 38 ;

 s413 =
  2500, 2495, 2490,
  2375, 2370, 2365,
  2250, 2245, 2240,
  2125, 2120, 2115 ;

 i414 =
  640000, 639980, 639960, 639940,
  632000, 631980, 631960, 631940,
  624000, 623980, 623960, 623940,
  616000, 615980, 615960, 615940 ;

 f421 =
  26244,
  26325,
  25515,
  25596,
  24786,
  24867,
  24057,
  24138 ;

 d422 =
  40000, 39990,
  40100, 40090,
  39000, 38990,
  39100, 39090,
  38000, 37990,
  38100, 38090,
  37000, 36990,
  37100, 37090 ;

 c423 =
  "@BD",
  "DFH",
  "HJL",
  "LNP",
  "PRT",
  "TVX",
  "XZ\\",
  "\\^`" ;

 b424 =
  64, 62, 60, 58,
  68, 66, 64, 62,
  56, 54, 52, 50,
  60, 58, 56, 54,
  48, 46, 44, 42,
  52, 50, 48, 46,
  40, 38, 36, 34,
  44, 42, 40, 38 ;

 s431 =
  2500,
  2525,
  2550,
  2375,
  2400,
  2425,
  2250,
  2275,
  2300,
  2125,
  2150,
  2175 ;

 i432 =
  640000, 639980,
  640400, 640380,
  640800, 640780,
  632000, 631980,
  632400, 632380,
  632800, 632780,
  624000, 623980,
  624400, 624380,
  624800, 624780,
  616000, 615980,
  616400, 616380,
  616800, 616780 ;

 f433 =
  26244, 26235, 26226,
  26325, 26316, 26307,
  26406, 26397, 26388,
  25515, 25506, 25497,
  25596, 25587, 25578,
  25677, 25668, 25659,
  24786, 24777, 24768,
  24867, 24858, 24849,
  24948, 24939, 24930,
  24057, 24048, 24039,
  24138, 24129, 24120,
  24219, 24210, 24201 ;

 d434 =
  40000, 39990, 39980, 39970,
  40100, 40090, 40080, 40070,
  40200, 40190, 40180, 40170,
  39000, 38990, 38980, 38970,
  39100, 39090, 39080, 39070,
  39200, 39190, 39180, 39170,
  38000, 37990, 37980, 37970,
  38100, 38090, 38080, 38070,
  38200, 38190, 38180, 38170,
  37000, 36990, 36980, 36970,
  37100, 37090, 37080, 37070,
  37200, 37190, 37180, 37170 ;

 c441 =
  "@",
  "D",
  "H",
  "L",
  "H",
  "L",
  "P",
  "T",
  "P",
  "T",
  "X",
  "\\",
  "X",
  "\\",
  "`",
  "d" ;

 b442 =
  64, 62,
  68, 66,
  72, 70,
  76, 74,
  56, 54,
  60, 58,
  64, 62,
  68, 66,
  48, 46,
  52, 50,
  56, 54,
  60, 58,
  40, 38,
  44, 42,
  48, 46,
  52, 50 ;

 s443 =
  2500, 2495, 2490,
  2525, 2520, 2515,
  2550, 2545, 2540,
  2575, 2570, 2565,
  2375, 2370, 2365,
  2400, 2395, 2390,
  2425, 2420, 2415,
  2450, 2445, 2440,
  2250, 2245, 2240,
  2275, 2270, 2265,
  2300, 2295, 2290,
  2325, 2320, 2315,
  2125, 2120, 2115,
  2150, 2145, 2140,
  2175, 2170, 2165,
  2200, 2195, 2190 ;

 i444 =
  640000, 639980, 639960, 639940,
  640400, 640380, 640360, 640340,
  640800, 640780, 640760, 640740,
  641200, 641180, 641160, 641140,
  632000, 631980, 631960, 631940,
  632400, 632380, 632360, 632340,
  632800, 632780, 632760, 632740,
  633200, 633180, 633160, 633140,
  624000, 623980, 623960, 623940,
  624400, 624380, 624360, 624340,
  624800, 624780, 624760, 624740,
  625200, 625180, 625160, 625140,
  616000, 615980, 615960, 615940,
  616400, 616380, 616360, 616340,
  616800, 616780, 616760, 616740,
  617200, 617180, 617160, 617140 ;
}
