netcdf bigr1 {
                // large last record variable
                // should work fine with classic format
                // should work fine with 64-bit offset format
dimensions:
	x = 100 ;
	y = 100 ;
	z = 100 ;
	t = UNLIMITED ;
variables:
	float x(x) ;
	float y(y) ;
	float z(z) ;
	float t(t) ;
	float var1(t) ;
	float var2(t, x, y, z) ;  // 4 GB OK since last record variable
data:
	var1 = 42 ;
}
