netcdf tst_charfill {
dimensions:
	STRING2 = 2 ;
	STRING4 = 4 ;
	STRING8 = 8 ;
	STRING16 = 16 ;
	STRING32 = 32 ;
	STRING256 = 256 ;
	iseq = UNLIMITED ; // (0 currently)
variables:
	int SEQUENCE(iseq) ;
		SEQUENCE:long_name = "PRG sequence number" ;
		SEQUENCE:units = "" ;
		SEQUENCE:conventions = "" ;
		SEQUENCE:_FillValue = 0 ;
		SEQUENCE:missing_value = 0 ;
		SEQUENCE:valid_min = 1 ;
		SEQUENCE:valid_max = 150000 ;
		SEQUENCE:tables = "results perform users comment" ;
	char IDENTIFIER(iseq, STRING32) ;
		IDENTIFIER:long_name = "Standard|sample identifier " ;
		IDENTIFIER:units = "" ;
		IDENTIFIER:conventions = "standard|G. species; left justified" ;
		IDENTIFIER:_FillValue = "";
		IDENTIFIER:tables = "results" ;

// global attributes:
		:version = "02a" ;
		:version_date = 20060501 ;
		:create_date = 20040323 ;
		:inew_start = 92586 ;
data:
 
SEQUENCE =
1
,2
,3
,4
,5
,6
,7
,8
,9
,10
,11
,12
,13
,14
,15
,16
,17
,18
,19
,20
,21
,22
,23
,24
,25
,26
,27
,28
,29
,30
,31
,32
,33
,34
,35
,36
;
}
