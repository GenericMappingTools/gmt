netcdf tst_group_data {
dimensions:
	dim = 4 ;
variables:
	float var(dim) ;
		var:units = "m/s" ;

// global attributes:
		:title = "for testing groups" ;
data:

 var = 1, 2, 3, 4 ;

group: g1 {
  dimensions:
  	dim = 1 ;
  variables:
  	float var(dim) ;
  		var:units = "km/hour" ;

  // group attributes:
  		:title = "in first group" ;
  data:

   var = 1 ;
  } // group g1

group: g2 {
  dimensions:
  	dim = 2 ;
  variables:
  	float var(dim) ;
  		var:units = "cm/sec" ;

  // group attributes:
  		:title = "in second group" ;
  data:

   var = 1, 2 ;

  group: g3 {
    dimensions:
    	dim = 3 ;
    variables:
    	float var(dim) ;
    		var:units = "mm/msec" ;
    	float var2(/dim, /g2/dim, dim) ;

    // group attributes:
    		:title = "in third group" ;
    data:

     var = 1, 2, 3 ;

     var2 =
  1, 2, 3,
  4, 5, 6,
  7, 8, 9,
  10, 11, 12,
  13, 14, 15,
  16, 17, 18,
  19, 20, 21,
  22, 23, 24 ;
    } // group g3
  } // group g2
}
