netcdf tst_comp {
types:
  compound obs_t {
    byte day ;
    short elev ;
    int count ;
    float relhum ;
    double time ;
    ubyte category ;
    ushort id ;
    uint particularity ;
    int64 attention_span ;
  }; // obs_t
dimensions:
	n = 3 ;
variables:
	obs_t obs(n) ;
		obs_t obs:_FillValue = {-99, -99, -99, -99, -99, 255, 65535, 4294967295, -9223372036854775806} ;
data:

 obs = {15, 2, 1, 0.5, 3600.01, 0, 0, 0, 0}, _, 
    {20, 6, 3, 0.75, 5000.01, 200, 64000, 4220002000, 9000000000000000000} ;
}
